library IEEE;
use ieee.std_logic_1164.all;